library ieee;
use ieee.std_logic_1164.all;

Entity processeur_monocycle_tb is
end entity;

Architecture TB of processeur_monocycle_tb is
  
  signal CLK, RST : std_logic;
  
  Begin
  
  process
    begin
    
      RST <= '1';
      clk <= '0';
      wait for 5 ns;
      RST <= '0';
      clk <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
      CLK <= '0';
      
      
      wait;
  end process;
  
  UUT: entity work.processeur_monocycle(RTL)  port map (CLK => CLK, RST => RST);
  
end TB;